
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
Use ieee.numeric_std.all;--displays a 6-bit unsigned value on the 7-segment displays.

Entity DispHex is
--code here

END DispHex ;

ARCHITECTURE operator OF DispHex IS
		--SIGNAL Sum : unsigned(7 downto 0);

Begin
--dispHEX accepts a 6-bit value, the 6 bits must be distributed between the two 7-segment decoders (Hint: use lab 3's segDecoder).

	--take sum here
	

END operator ;
